module top(
  );

  initial
  begin
    $dumpfile("ipc.vcd");
    $dumpvars(1,top);
  end


endmodule
