module top(
  );
 
  
endmodule