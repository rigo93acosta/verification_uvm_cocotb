module top(
  );

  initial
  begin
    $dumpfile("classIPC.vcd");
    $dumpvars(1,top);
  end


endmodule
